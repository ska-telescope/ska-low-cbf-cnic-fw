--------------------------------------------------------------------------------
--
--  This file was automatically generated using ARGS config file <lib>.peripheral.yaml
--
--
--
--
--------------------------------------------------------------------------------

library ieee, axi4_lib, common_lib;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use axi4_lib.axi4_lite_pkg.ALL;
use common_lib.common_pkg.ALL;

-------------------------------------------------------------------------------
package <lib_name>_reg_pkg is

   ---------------------------------------------------------------------------
   --                        COMPONENT DECLARATIONS                         --
   ---------------------------------------------------------------------------



    ---------------------------------------------------------------------------
    --                CONSTANT, TYPE AND GENERIC DEFINITIONS                 --
    ---------------------------------------------------------------------------


    <{constant_statements}>

    <{type_statements}>

end <lib_name>_reg_pkg;

-------------------------------------------------------------------------------
package body <lib_name>_reg_pkg is


   ---------------------------------------------------------------------------
   --                 FUNCTION/PROCEDURE DEFINITIONS                        --
   ---------------------------------------------------------------------------


end <lib_name>_reg_pkg;
-------------------------------------------------------------------------------



